module main

fn main() {
	mut strings := ['hello', 'world']
	for idx, el in strings {
		println('${idx} ${el}')
		println('${idx} ${strings[idx]}')
	}
	for idx, _ in strings {
		println(idx)
	}
	for _ in strings {
		println('hello')
	}
	for i, _ in [2]int{} {
		for j, _ in [2]int{} {
			println('hello2')
		}
	}
}
