module main

fn main() {
	mut a := 1 & ~2
	mut b := 1 + 2 + 3 + -4
}
