module main

fn main() {
	println('Hello World')
	mut ok := Test1{}
	ok.a.test()
	println('okkk')
}

struct Test1 {
pub mut:
	a Test2
}

struct Test2 {
}

fn (t Test2) test() {
	println('Test')
}
