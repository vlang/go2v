module main

fn main() {
	func()
}

fn func() {
}
