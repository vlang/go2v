module main

fn main() {
	if true {
		println('true')
	} else {
		println(2 + 3)
	}
}
